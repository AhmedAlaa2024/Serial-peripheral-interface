module Master(CS, SCLK, MOSI, MISO);


endmodule
