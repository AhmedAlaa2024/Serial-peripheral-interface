module Slave_TB();



endmodule