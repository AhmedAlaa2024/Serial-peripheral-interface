module Slave(CS, SCLK, SDI, SDO);



endmodule