module Master_TB();


endmodule