module Slave(
	reset,
	slaveDataToSend, slaveDataReceived,
	SCLK, CS, MOSI, MISO
);



endmodule